`timescale 1ns / 1ps

module PS2MOUSE(CLK,RST,PS2CLK,PS2DATA,STREAM,FAIL,DatoRec);
	input CLK,RST;
	inout PS2CLK,PS2DATA;
	output wire STREAM,FAIL;
	output wire [7:0] DatoRec;

//Redes
	wire PS2CLKO,PS2DATAO;
	wire ENABC,ENABD;
	Buffer1bit BCLK(PS2CLKO,ENABC,PS2CLK);
	Buffer1bit BDATA(PS2DATAO,ENABD,PS2DATA);
	
	wire PS2CLKR,PS2CLKE,PS2DATAR,PS2DATAE;
	wire ENABCR,ENABCE,ENABDR,ENABDE;
	
	assign PS2CLKO=PS2CLKR&PS2CLKE;
	assign PS2DATAO=PS2DATAR&PS2DATAE;
	assign ENABC=ENABCR|ENABCE;
	assign ENABD=ENABDR|ENABDE;
	
//FSM de recepcion
	FSMPS2MOUSE FSMREC(CLK,RST,PS2CLK,PS2DATA,PS2CLKR,PS2DATAR,DatoRec,STREAM,FAIL,ENABCR,ENABDR);

//FSM de ENVIO
	FSMPS2MOUSE2 FSMENV(CLK,RST,STREAM,PS2CLKE,PS2DATAE,ENABCE,ENABDE);
	
endmodule
