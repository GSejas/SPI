`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
module FSMControlPS2(
    input ena,
	 input rst,
	 input clk,
    output data);
//Declaracion de las entradas



