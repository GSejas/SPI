`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
module PS2_Rx(clk, rst, fall_edge,ps2_d, rx_done,  DataOut);


endmodule
